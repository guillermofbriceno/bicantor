module execute
(
    input wire [31:0]        inst0_i,
    input wire [31:0]        inst1_i,
    input wire [`CTRL_BUS]   ctrl0_i,
    input wire [`CTRL_BUS]   ctrl1_i,
    input wire [31:0]        rs1_data0_i,
    input wire [31:0]        rs2_data0_i,
    input wire [31:0]        rs1_data1_i,
    input wire [31:0]        rs2_data1_i
     
);

 endmodule
