module lsu
(
    input [31:0] alu0_out_i,
    input [31:0] alu1_out_i
);

endmodule
